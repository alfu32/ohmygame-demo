module ohmygame

fn test_drawing_context_2d_create(){
	vp:=drawing_context_2d_create(120,40," ")

	dump(vp)
}

