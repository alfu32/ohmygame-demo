module main

// import ohmygame

pub fn make_player_ship(){}