module ohmygame


pub fn test_pad_end() {
	a:="abcd"
	b:=pad_end(a,3,">")
}
pub fn test_pad_start() {
	a:="abcd"
	b:=pad_start(a,3,">")
}